module DebounceTest;


/*[TestModule --module Debounce]*/


initial begin

    #5000;


    /*[PressButton]*/

    /*[PressButton]*/

    /*[PressButton]*/

    /*[PressButton]*/

    /*[PressButton]*/

    /*[PressButton]*/

    /*[PressButton]*/

    #50000;
    $finish;
    
end
endmodule